LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;

ENTITY NIOSII IS
    PORT (
        -- 50 MHz clock to drive out system
        CLOCK_50 : IN STD_LOGIC;
        -- Array of 8 green LEDs on the development board for output
        LEDG : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
END NIOSII;

ARCHITECTURE Structure OF NIOSII IS
    -- Design ports to interact with the generated architecture
    COMPONENT NIOSII_DE2
        PORT (
            clk_50 : IN STD_LOGIC;
            reset_n : IN STD_LOGIC;
            out_port_from_the_pio_led : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
        );
    END COMPONENT;

BEGIN
--Instantiate the Nios II system entity generated by the SOPC Builder
    Def: NIOSII_DE2 PORT MAP (CLOCK_50, '1', LEDG);

END Structure;
